module Icache
(
    input clk,
    input rst,

    input icache_valid,
    input [63:0] inst_in_data_32,
    input [16*32-1:0] inst_in_data_shortcut,
    input [31:0] inst_addr,
    input inst_en,
    //input data_in_ready,
    input mem_stop,
    input dcache_busy,
    input icache_ready,
    input read_shortcut,
    output [31:0] inst_read_addr,
    output inst_read_req,
    output reg [31:0] inst_out_data
);

wire [15:0]hit;
reg [25:0] tag [15:0]   ;         //total 16 index  therefore ,22 bits tag
reg [511:0] inst_store [15:0];   //16 is a set
reg [9:0] offset;
wire [9:0] offset_wire;
reg [31:0] inst_addr_pre;
wire [31:0] inst_addr_sel;
assign inst_addr_sel = icache_state == 2'd1 |mem_stop ?inst_addr_pre : inst_addr;
//generated by script
assign hit[0] = tag[0] == inst_addr_sel[31:6];
assign hit[1] = tag[1] == inst_addr_sel[31:6];
assign hit[2] = tag[2] == inst_addr_sel[31:6];
assign hit[3] = tag[3] == inst_addr_sel[31:6];
assign hit[4] = tag[4] == inst_addr_sel[31:6];
assign hit[5] = tag[5] == inst_addr_sel[31:6];
assign hit[6] = tag[6] == inst_addr_sel[31:6];
assign hit[7] = tag[7] == inst_addr_sel[31:6];
assign hit[8] = tag[8] == inst_addr_sel[31:6];
assign hit[9] = tag[9] == inst_addr_sel[31:6];
assign hit[10] = tag[10] == inst_addr_sel[31:6];
assign hit[11] = tag[11] == inst_addr_sel[31:6];
assign hit[12] = tag[12] == inst_addr_sel[31:6];
assign hit[13] = tag[13] == inst_addr_sel[31:6];
assign hit[14] = tag[14] == inst_addr_sel[31:6];
assign hit[15] = tag[15] == inst_addr_sel[31:6];

assign inst_read_req = (hit==16'd0) && inst_en;
assign inst_read_addr = {inst_addr_sel[31:6],6'd0};

//The following is the replacement algorithm
reg [3:0] replace_index;
always @(posedge clk)
begin
    if(rst) begin
        replace_index <= 4'd0;
    end
    else begin
        //$display("%d\n",inst_addr_sel);
        replace_index <= replace_index +4'd1;   
    end
        
end
wire [3:0] hit_index;
find_index find_index_hit(
    .data(hit),
    .index(hit_index)
);
reg [1:0] icache_state;
reg [3:0] index_replace_real;
reg [3:0] index_in;
reg [3:0] replace_index_reg ;
always @(posedge clk) begin
    if(rst) begin
        for(int i=0;i<16;i++) begin
            inst_store[i] <=512'd0;
        end
        for(int j=0;j<16;j++) begin
            tag[j] <= 26'd0;
        end
        icache_state <= 2'd0;
        inst_addr_pre <= 32'd0;
    end
    else if(icache_state == 2'd1 && icache_valid) begin
        inst_store[replace_index_reg][({2'd0,index_in}+6'd1)*32-1-:32] <= index_in[0] == 0?inst_in_data_32[31:0]:inst_in_data_32[63:32];
        index_in <= index_in +1;
        if(icache_ready) begin
            icache_state <= 2'd0;
            tag[replace_index_reg] <= inst_addr_sel[31:6];
        end
        if(inst_addr_sel[5:2] == index_in) begin
            inst_out_data <= index_in[0] == 0?inst_in_data_32[31:0]:inst_in_data_32[63:32];
        end
        
    end
    else if(dcache_busy)begin 
    end
    else if(icache_state == 2'd0) begin //ready state
        if(inst_read_req && ~read_shortcut)begin   //there should be a not busy
            icache_state <= 2'd1; // wait state
            inst_addr_pre <= inst_addr;
            index_in <= 4'd0;
            replace_index_reg <= replace_index;
        end
        else if(inst_read_req && read_shortcut) begin
            inst_out_data <= inst_in_data_shortcut[offset_wire-1-:32];
            inst_store[replace_index] <= inst_in_data_shortcut;
            tag[replace_index] <= inst_addr_sel[31:6];
            inst_addr_pre <= inst_addr;
        end
        else begin
            inst_out_data <= inst_store[hit_index][offset_wire-1-:32];
            inst_addr_pre <= inst_addr;
        end
    end
end
assign offset_wire = ({6'd0,{inst_addr_sel[5:2]}}+10'd1) <<5;


endmodule