module mul_32 (
    input [31:0] src1,
    input [31:0] src2,

    output [63:0] output1
);
    assign output1 = ({32'd0,(src1[0] ? src2 : 32'd0)} << 0) +
                    ({32'd0,(src1[1] ? src2 : 32'd0)} << 1) +
                    ({32'd0,(src1[2] ? src2 : 32'd0)} << 2) +
                    ({32'd0,(src1[3] ? src2 : 32'd0)} << 3) +
                    ({32'd0,(src1[4] ? src2 : 32'd0)} << 4) +
                    ({32'd0,(src1[5] ? src2 : 32'd0)} << 5) +
                    ({32'd0,(src1[6] ? src2 : 32'd0)} << 6) +
                    ({32'd0,(src1[7] ? src2 : 32'd0)} << 7) +
                    ({32'd0,(src1[8] ? src2 : 32'd0)} << 8) +
                    ({32'd0,(src1[9] ? src2 : 32'd0)} << 9) +
                    ({32'd0,(src1[10] ? src2 : 32'd0)} << 10) +
                    ({32'd0,(src1[11] ? src2 : 32'd0)} << 11) +
                    ({32'd0,(src1[12] ? src2 : 32'd0)} << 12) +
                    ({32'd0,(src1[13] ? src2 : 32'd0)} << 13) +
                    ({32'd0,(src1[14] ? src2 : 32'd0)} << 14) +
                    ({32'd0,(src1[15] ? src2 : 32'd0)} << 15) +
                    ({32'd0,(src1[16] ? src2 : 32'd0)} << 16) +
                    ({32'd0,(src1[17] ? src2 : 32'd0)} << 17) +
                    ({32'd0,(src1[18] ? src2 : 32'd0)} << 18) +
                    ({32'd0,(src1[19] ? src2 : 32'd0)} << 19) +
                    ({32'd0,(src1[20] ? src2 : 32'd0)} << 20) +
                    ({32'd0,(src1[21] ? src2 : 32'd0)} << 21) +
                    ({32'd0,(src1[22] ? src2 : 32'd0)} << 22) +
                    ({32'd0,(src1[23] ? src2 : 32'd0)} << 23) +
                    ({32'd0,(src1[24] ? src2 : 32'd0)} << 24) +
                    ({32'd0,(src1[25] ? src2 : 32'd0)} << 25) +
                    ({32'd0,(src1[26] ? src2 : 32'd0)} << 26) +
                    ({32'd0,(src1[27] ? src2 : 32'd0)} << 27) +
                    ({32'd0,(src1[28] ? src2 : 32'd0)} << 28) +
                    ({32'd0,(src1[29] ? src2 : 32'd0)} << 29) +
                    ({32'd0,(src1[30] ? src2 : 32'd0)} << 30) +
                    ({32'd0,(src1[31] ? src2 : 32'd0)} << 31) ;
endmodule