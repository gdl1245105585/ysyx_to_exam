module AXI4 (


    
);
    
assign AWPROT = 3'b011;
endmodule